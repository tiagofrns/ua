library IEEE;
use IEEE.STD_LOGIC_1164;

entity ShiftRegister4 in
	port(			
		clk: in std_logic;
		sin: in std_logic;
		dataOut: out std_logic_vector(3 downto 0)
	
	);
	
end ShiftRegister4;



architecture Shell of ShiftRegister4 is

begin






end Shell;